library ieee;
use ieee.std_logic_1164.all;

--! Used data types for MCU
package data_types is

	constant signal R0 : std_logic_vector := 0;
	constant signal R1 : std_logic_vector := 1;
	constant signal R2 : std_logic_vector := 2;
	constant signal R3 : std_logic_vector := 3;
	

end package;
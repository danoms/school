package basic_bit_blocks is

	


end package;